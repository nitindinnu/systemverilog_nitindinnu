module name(
    port_list
);
    
endmodule