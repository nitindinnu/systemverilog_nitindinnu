module dynamic_array_test(
);
/*create a 32x32 bit memoryusing dynamic array & fill memory with your own data & read then extend it to 32x64 memory .check whether old data is there or not*/
    bit [31:0]dynamicarray[];

    initial begin
        dynamicarray=new[32];
        foreach (dynamicarray[i]) begin
            dynamicarray[i]=$random;
        end
        $display("elements of 32 %p",dynamicarray);
        dynamicarray=new[64](dynamicarray);
        $display("elements of 64 %p",dynamicarray);
/*
# Loading work.dynamic_array_test(fast)

# elements of 32 '{303379748, 3230228097, 2223298057, 2985317987, 112818957, 1189058957, 2999092325, 
2302104082, 15983361, 114806029, 992211318, 512609597, 
1993627629, 1177417612, 2097015289, 3812041926, 3807872197, 3574846122, 1924134885, 
3151131255, 2301810194, 1206705039, 2033215986, 3883308750, 4093672168, 3804909253, 777537884, 3733858493, 2527811629, 
2997298789, 2985255523, 91457290}

# elements of 64 '{303379748, 3230228097, 2223298057, 2985317987, 112818957, 1189058957, 2999092325, 2302104082, 15983361, 114806029,
 992211318, 512609597, 1993627629, 1177417612, 2097015289, 3812041926, 3807872197, 3574846122, 1924134885, 
3151131255, 2301810194, 1206705039, 2033215986, 3883308750, 4093672168, 3804909253, 777537884, 3733858493,
 2527811629, 2997298789, 2985255523, 91457290, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
0, 0, 0, 0,0, 0, 0, 0, 0, 0}
*/

    end
endmodule