module store_array_in_queue(
);
    /*Ex : `arr[8] = '{5,6,8,3,4,9,7,2}'` is the input sort & store in the queue `Q1[$]` and display that queue*/

    reg[2:0] arr;
endmodule