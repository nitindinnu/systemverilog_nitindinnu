module (
    port_list
);
    
endmodule