class generator;
    
endclass