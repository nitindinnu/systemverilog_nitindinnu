//  Module: 02tasks
//
module tasks01 ();//! static task

    
endmodule: tasks01


module task02();//! automatic task
    
endmodule

module task03();//! global task
    
endmodule

module task04(); //! disable task
    
endmodule
